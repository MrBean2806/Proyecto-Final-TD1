library verilog;
use verilog.vl_types.all;
entity Filtro_Rebote_tb is
end Filtro_Rebote_tb;
