library verilog;
use verilog.vl_types.all;
entity Drv_display_tb is
end Drv_display_tb;
